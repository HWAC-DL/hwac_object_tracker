
`timescale 1ns / 1ps

module shift_reg
    (
        clk,

        enable,
        data_in,
        data_out
    );

//-------------------------------------------------------------------------------------------------
// Global constant headers
//-------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
// Parameter definitions
//-------------------------------------------------------------------------------------------------
    parameter                                                   CLOCK_CYCLES = 8;
    parameter                                                   DATA_WIDTH   = 128;
//-------------------------------------------------------------------------------------------------
// Localparam definitions
//-------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
// I/O signals
//-------------------------------------------------------------------------------------------------
    input                                                       clk;

    input                                                       enable;
    input       [DATA_WIDTH-1:0]                                data_in;
    output 		[DATA_WIDTH-1:0]                                data_out;
//-------------------------------------------------------------------------------------------------
// Internal wires and registers
//-------------------------------------------------------------------------------------------------
    reg         [CLOCK_CYCLES-1:0]                              shift_reg [DATA_WIDTH-1:0];
//-------------------------------------------------------------------------------------------------
// Implementation
//-------------------------------------------------------------------------------------------------

   genvar i;
   generate
        for (i=0; i < DATA_WIDTH; i=i+1) begin: shift_blk
            always @(posedge clk) begin
                if(enable) begin
                    shift_reg[i] <= {shift_reg[i][CLOCK_CYCLES-2:0], data_in[i]};
                end
            end
            assign data_out[i] = shift_reg[i][CLOCK_CYCLES-1];
        end
   endgenerate

endmodule