`timescale 1ns / 1ps

module vector2index
    (
        vector_in,
        index_out,
        contains_valid_index_out
    );

//-------------------------------------------------------------------------------------------------
// Global constant headers
//-------------------------------------------------------------------------------------------------
    `include "util_funcs.v"
//-------------------------------------------------------------------------------------------------
// Parameter definitions
//-------------------------------------------------------------------------------------------------
    parameter   VECTOR_WIDTH    = 8;
//-------------------------------------------------------------------------------------------------
// Localparam definitions
//-------------------------------------------------------------------------------------------------
    localparam  INDEX_WIDTH     = count2width(VECTOR_WIDTH);
//-------------------------------------------------------------------------------------------------
// I/O signals
//-------------------------------------------------------------------------------------------------
    input       [VECTOR_WIDTH-1:0]  vector_in;
    output reg  [INDEX_WIDTH-1:0]   index_out;      //syntheized to a wire not a reg
    output reg                      contains_valid_index_out;
//-------------------------------------------------------------------------------------------------
// Internal wires and registers
//-------------------------------------------------------------------------------------------------
    integer                     i;
//-------------------------------------------------------------------------------------------------
// Implementation
//-------------------------------------------------------------------------------------------------
    always@(*) begin
        index_out = {INDEX_WIDTH{1'b0}};
        contains_valid_index_out    = (|vector_in) ? 1'b1 : 1'b0;
        for (i=(VECTOR_WIDTH-1); i>=0; i=i-1) begin
            if (vector_in[i] == 1'b1) begin
                index_out = i;
            end
        end
    end

endmodule
